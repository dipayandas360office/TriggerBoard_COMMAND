library IEEE;
library UNISIM;
use UNISIM.VComponents.all;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity Trigger is 
    generic (
        baud                : positive := 921600;
        clock_frequency     : positive := 100_000_000
    );
port (
--    clock : in std_logic;
    clk_in                  : in std_logic;
    clk_out                 : out std_logic;
    trig_in                 : in std_logic;
    trig_out1               : out std_logic;
    trig_out2               : out std_logic;
    bin_number              : in std_logic_vector (3 downto 0);
    usb_rs232_rxd           : in      std_logic;
    usb_rs232_txd           : out     std_logic;
    reset_in                : in std_logic;
    led_signal              : out std_logic
);
end Trigger;

architecture behav of Trigger is 
signal clk_40 , clk_100 , clk_400 : std_logic:='0';
signal reset_s : std_logic :='0';
signal mono_out : std_logic := '0' ;
signal mono_on : std_logic := '0';
signal count : integer := 0;
signal trig_out : std_logic := '0';
signal clk_locked : std_logic;
signal trig_in_d1 , trig_in_d2 , trig_rise , clk_in_d1 , clk_in_d2 , clk_in_rise ,trig_out_and: std_logic := '0';
signal count_bin    : unsigned(3 downto 0):="0000";
signal trig_out_buf ,gate : std_logic;

    -----Rx Tx of USB--------------------------------------------------------------------------------------
signal tx, rx, rx_sync, reset, reset_sync       : std_logic;
signal fifo_data_in_stb_t , fifo_data_out_stb   : std_logic;
signal  fifo_data_in_t,fifo_data_out,command    : std_logic_vector ( 7 downto 0);
signal fifo_empty, fifo_full_t                  : std_logic;
signal sendLogic , command_execute               : std_logic := '0';

    -- Component declaration for clk_wiz_0
component clk_wiz_0
    port(
       clk_out1   : out std_logic;
       clk_out2   : out std_logic;
       reset      : in  std_logic;
       locked     : out std_logic;
       clk_in1    : in std_logic
    );
end component;

    component UartCommand is
    generic (
        baud                : positive;
        clock_frequency     : positive
    );
    port(  
    clock                   : in   std_logic;
    reset                   : in   std_logic;  
    rx                      : in   std_logic;
    tx                      : out  std_logic;
    fifo_empty              : out  std_logic;
    fifo_full_t             : out  std_logic;
    fifo_data_in_stb_t      : in   std_logic;
    fifo_data_out_stb       : in   std_logic;
    fifo_data_in_t          : in   std_logic_vector(7 downto 0);
    fifo_data_out           : out  std_logic_vector(7 downto 0)
    );
end component UartCommand;
 
begin

    ----------------------------------------------------------------------------
--  USB Uart_Command instantiation
----------------------------------------------------------------------------
UartCommandInstance : UartCommand
generic map (
    baud                => baud,
    clock_frequency     => clock_frequency
)
port map (  
    clock               => clk_100,
    reset               => reset,    
    rx                  => rx,
    tx                  => tx,
    fifo_empty          => fifo_empty,
    fifo_full_t         => fifo_full_t,
    fifo_data_in_stb_t  => fifo_data_in_stb_t,
    fifo_data_out_stb   => fifo_data_out_stb,
    fifo_data_in_t      => fifo_data_in_t ,   
    fifo_data_out       => fifo_data_out
   
);

    ClockGen : clk_wiz_0
    port map(
        clk_out1  => clk_400,
        clk_out2  => clk_100,
        reset     => reset_s,
        clk_in1   => clk_in,
        locked    => clk_locked
    );

    OBUF_inst : OBUF
        generic map (
            DRIVE => 12,
            IOSTANDARD => "LVCMOS33",
            SLEW => "FAST"
        )
        port map(
            I => clk_in,
            O => clk_out
        );

trig    : process (clk_400) 
          begin
          if rising_edge(clk_400) then
              if (reset_s ='1') then
                    count_bin <= "0000";
--                    count <= 0;
--                    mono_on    <= '0';
--                    trig_out   <= '0';
              else
                  if count_bin = 9 then
                     count_bin <= "0000";
                  else 
                    count_bin <= count_bin +1; 
                  end if;
                  
                  trig_in_d1 <= trig_in;
                  trig_in_d2 <= trig_in_d1;
                  
--                  clk_in_d1 <= clk_in;
--                  clk_in_d2 <= clk_in_d1;
                                                      
--                  if (count_bin >= "0011" and count_bin <="0100"  ) then ------------- select the bin (phase)
                 if (bin_number = "1111") then 
                    gate <= '1';
                 else                                     
                      if (count_bin = unsigned(bin_number)) then ------------- select the bin (phase)
                        gate <='1';
                      else
                        gate <= '0';
                      end if;
                 end if; 
               end if;
          end if;
       end process; 
        
monoshot : process (clk_400)
       begin
           if rising_edge(clk_400) then
               if (reset_s = '1') then
                   count <= 0;
                   trig_out_buf <= '0';
--               elsif (gate = '1' and trig_rise = '1') then
               elsif (gate = '1' and trig_in = '1') then -- ANDed with Trig_in
                   count <= 0;
                   trig_out_buf <= '1';
               elsif (trig_out_buf = '1') then
                   if (count < 39) then
                       count <= count + 1;
                   else
                       count <= 0;
                       trig_out_buf <= '0';
                   end if;
               end if;
           end if;
       end process;

    ----------------------------------------------------------------------------
       -- Deglitch inputs
       ----------------------------------------------------------------------------
deglitch : process (clk_100)
begin
   if rising_edge(clk_100) then
       rx_sync         <= usb_rs232_rxd;
       rx              <= rx_sync;
       reset_sync      <= reset_in;
       reset           <= reset_sync;
       usb_rs232_txd   <= tx;
   end if;
end process;

Loopbak : process(clk_100)
begin
    if rising_edge(clk_100) then
         ----------------------Reset logic -------------------------------------   
            if reset = '1' then
                fifo_data_out_stb       <= '0';
                fifo_data_in_stb_t      <= '0';  
     -------------------------------------------------------------------------
            else
          -----------Transmit and receive  initialize 
                fifo_data_out_stb       <= '0';
                fifo_data_in_stb_t      <= '0';
                
---------------Loop back code -----------------------------                
                 if fifo_EMPTY = '0' then
                     if sendlogic = '0' then
                         fifo_data_out_stb <= '1';
                         command   <= fifo_data_out;
                         sendlogic <= sendlogic xor '1';
                     elsif sendlogic = '1' then
                        if fifo_full_t = '0' then
                            fifo_data_in_stb_t <= '1';
                            fifo_data_in_t     <= command;
                            sendlogic <= sendlogic xor '1';
                        end if;
                     end if;
                 end if;
------------------------Loop back code ends -----------------
                 ---------------------------Reading the Command--------------------------------------------------
                if fifo_empty = '0' and sendLogic = '0' then
                    fifo_data_out_stb <= '1';
                
                    -- Simple command (like 0x31 or 0x32)
                    if (fifo_data_out = x"31" or fifo_data_out = x"32") and HVDB_cmd_on = "00" then
                        command_execute <= '1';
                        command <= fifo_data_out;
                        sendLogic <= sendLogic xor '1';  
                    -- First byte of HVDB command (ignored)
                    elsif fifo_data_out = x"61" or fifo_data_out = x"62" then
                        HVDB_cmd_on <= "01";  -- move to next byte
                        sendLogic <= sendLogic xor '1';  
                        command_HVDB(31 downto 24) <= fifo_data_out;
                    -- Second byte of HVDB command (first useful byte)
                    elsif HVDB_cmd_on = "01" then
                        command_HVDB(23 downto 16) <= fifo_data_out;  -- store as high byte
                        HVDB_cmd_on <= "10";                           -- reset FSM
                        sendLogic <= sendLogic xor '1';    
                    -- Third byte of HVDB command (second useful byte)
                    elsif HVDB_cmd_on = "10" then
                        command_HVDB(15 downto 8) <= fifo_data_out;   -- store as low byte            
                        HVDB_cmd_on <= "11";                           -- reset FSM
                        sendLogic <= sendLogic xor '1';               -- signal complete    
                    -- Fourth byte of HVDB command (third useful byte)
                    elsif HVDB_cmd_on = "11" then
                        command_HVDB(7 downto 0) <= fifo_data_out;   -- store as low byte
                        HVDB_control_in_s <= '1';                     -- trigger processing
                        HVDB_cmd_on <= "00";                           -- reset FSM
                        sendLogic <= sendLogic xor '1';               -- signal complete
                    
                
                    else
                        command_execute <= '0';
                        sendLogic <= sendLogic xor '1';
                        if fifo_data_out = x"33" then
                            resetTimer <= '1';
                        end if;
                    end if;
                                        
                 elsif fifo_empty_r_ethernet = '0' and sendLogic = '0'  then
                    fifo_data_out_stb_r_ethernet       <= '1';
                    if fifo_data_out_r_ethernet = x"31" or fifo_data_out_r_ethernet = x"32" then
                        command_execute <= '1';
                        command <= fifo_data_out_r_ethernet;
                    else    
                        command_execute <= '0';
                        sendLogic <= sendLogic xor '1';
                        if fifo_data_out_r_ethernet = x"33" then
                        resetTimer <= '1';
                        end if;
                    end if;
                elsif sendLogic = '1' then
                    sendLogic <= sendLogic xor '1';
                end if;
              end if;
             end if;
    end process;
             end if;
    end if;
end process;    

command_exec : process( clk_100)
begin
    if rising_edge(clk_100) then 
        if (command = x"31" ) then
            led_signal <= '1';
        elsif command = x"32" then
            led_signal <= '0';
        end if;
    end if;

end process;

--trig_out1 <= gate;
trig_out1 <= trig_out_buf;                   
reset_s <= reset_in;   
trig_rise <= trig_in_d1 and not trig_in_d2;   -- rising edge detect  
trig_out_and <= gate and trig_rise;
clk_40 <= clk_in;
--trig_out2 <= trig_out_and;
trig_out2 <= trig_out_buf;
--clk_out <= clk_40;
--counterOut <= std_logic(count_bin(2));
end behav;
